module gate(a, b, y);
input a;
output y;
assign y = ~a;
endmodule
